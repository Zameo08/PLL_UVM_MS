//------------------------------------------------------------------------------
//
// registers transaction enums, parameters, and events
//
//------------------------------------------------------------------------------

// enum to control coverage
typedef enum bit {COV_ENABLE, COV_DISABLE} cover_e;
