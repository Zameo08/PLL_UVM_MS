package pll_pkg;

  import uvm_pkg::*;
  import uvm_ms_pkg::*;
  `include "uvm_macros.svh"

  `include "pll_types.sv"
  `include "pll_transaction.sv"
  `include "pll_ms_transaction.sv"
  `include "pll_bridge_proxy.sv"
  `include "pll_sequencer.sv"
  `include "pll_monitor.sv"
  `include "pll_ms_source_monitor.sv"
  `include "pll_driver.sv"
  `include "pll_ms_source_driver.sv"
  `include "pll_base_seq.sv"
  `include "pll_base_ms_seq.sv"
  `include "pll_nested_seq.sv"
  `include "pll_ms_source_transaction_seq.sv"
  `include "pll_ms_source_nested_seq.sv"
  `include "pll_agent.sv"
  `include "pll_env.sv"

endpackage : pll_pkg