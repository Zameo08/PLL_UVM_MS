//------------------------------------------------------------------------------
//
// osc_ms transaction enums, parameters, and events
//
//------------------------------------------------------------------------------

typedef enum bit {OSC_MS_DRIVE, OSC_MS_SAMPLE } osc_ms_data_type_e;
